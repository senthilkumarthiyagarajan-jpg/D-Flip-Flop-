.title KiCad schematic
ID_in_plt1 D_IN PLOT 1
VDIN1 D_IN GND pulse(0 5 0 1ns 1ns 20ns 40ns)
M2N1 Net-_M1N1-Pad3_ D_IN GND GND eSim_MOS_N
VCLKIN1 /CLK GND pulse(0 5 0 1n 1n 5n 10n)
M1N1 QBAR_OUT /CLK Net-_M1N1-Pad3_ GND eSim_MOS_N
CLKINPLT1 /CLK PLOT 3
M3N1 Q_OUT QBAR_OUT GND GND eSim_MOS_N
M5N1 Net-_M4N1-Pad3_ Q_OUT GND GND eSim_MOS_N
out_bar1 QBAR_OUT PLOT5
M4N1 QBAR_OUT /CLKB Net-_M4N1-Pad3_ GND eSim_MOS_N
M2P1 Net-_M1P1-Pad3_ /CLKB QBAR_OUT /VDD eSim_MOS_P
M1P1 /VDD D_IN Net-_M1P1-Pad3_ /VDD eSim_MOS_P
CLKBINPLT1 /CLKB PLOT2
VCLKBIN1 /CLKB GND pulse(5 0 0 1n 1n 5n 10n)
M3P1 /VDD QBAR_OUT Q_OUT /VDD eSim_MOS_P
M4P1 /VDD Q_OUT Net-_M4P1-Pad3_ /VDD eSim_MOS_P
out1 Q_OUT PLOT4
M5P1 Net-_M4P1-Pad3_ /CLK QBAR_OUT /VDD eSim_MOS_P
VDD1 /VDD GND dc 5
.end
